`define TEST_COUNT 14
`define TRACE_FILE_PATH "./lab2.data/lab2_cpu_trace"
`define INST_FILE_PATH  "./lab2.data/lab2_inst_data"
`define DATA_FILE_PATH  "./lab2.data/lab2_data_data"
`define GPRS_FILE_PATH  "./lab2.data/lab2_reg_data"
